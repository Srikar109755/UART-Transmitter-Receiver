`timescale 1ns / 1ps


`include "Baud_Gen.sv"
`include "UART_TX.sv"
`include "UART_RX.sv"